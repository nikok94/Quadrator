IntToFloat_inst : IntToFloat PORT MAP (
		clock	 => clock_sig,
		dataa	 => dataa_sig,
		result	 => result_sig
	);
